// Control unit - Signed, 9662e103-129a

module cu ();

endmodule