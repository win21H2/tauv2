// Interface - Signed, 9662e103-129a

module interface ();

endmodule