// Arithmetic logic unit - Signed, 9662e103-129a

module alu ();

endmodule