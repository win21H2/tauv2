// Program counter - Signed, 9662e103-129a

module pc ();

endmodule