// Register file - Signed, 9662e103-129a

module rf ();

endmodule